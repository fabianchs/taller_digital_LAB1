module tb_full_adder_mega_extended;

    logic[63:0] A,B;
    logic Cin;
    logic Cout;
    logic [63:0]S;
    
    full_adder_mega_extended dut(
    
    .A (A),
    .B (B),
    .Cin (Cin),
    .Cout (Cout),
    .S (S)
    
    );
    
    initial begin
        
        A<=64'b0010100100101001001010010010100100101001001010010010100100101001;
        B<=64'b0010110100101101001011010010110100101101001011010010110100101101;
        Cin<=0;
        #10
        A<=64'b0110100101101001011010010110100101101001011010010110100101101001;
        B<=64'b1010110110101101101011011010110110101101101011011010110110101101;
        Cin<=1;
        #10
        A<=64'b1110111111101111111011111110111111101111111011111110111111101111;
        B<=64'b1010011110100111101001111010011110100111101001111010011110100111;
        Cin<=1;
        #10
        A<=64'b0111110101111101011111010111110101111101011111010111110101111101;
        B<=64'b1010110110101101101011011010110110101101101011011010110110101101;
        Cin<=0;
        #10
        A<=64'b0100110101001101010011010100110101001101010011010100110101001101;
        B<=64'b0110110101101101011011010110110101101101011011010110110101101101;
        Cin<=0;
        #10
        A<=64'b0111010101110101011101010111010101110101011101010111010101110101;
        B<=64'b1110010111100101111001011110010111100101111001011110010111100101;
        Cin<=0;
        #10
        A<=64'b0100110101001101010011010100110101001101010011010100110101001101;
        B<=64'b1011110110111101101111011011110110111101101111011011110110111101;
        Cin<=0;
        #10
        $finish;
    
    end
    
endmodule