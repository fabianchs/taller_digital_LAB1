`timescale 1ns / 1ps


module tb_mux_4_1;

    logic [15:0]in0;
    logic [15:0]in1;
    logic [15:0]in2;
    logic [15:0]in3;
    logic [1:0]sel;
    logic [15:0] out;


    mux_4_1 dut(
    
    .in0 (in0),
    .in1 (in1),
    .in2 (in2),
    .in3 (in3),
    .sel (sel),
    .out (out));
    
    initial begin 
        in0<=1;
        in1<=1;
        in2<=1;
        in3<=1;
        sel<=0;
        #10
        in0<=1;
        in1<=0;
        in2<=1;
        in3<=0;
        sel<=1;
        #10
        in0<=0;
        in1<=1;
        in2<=1;
        in3<=1;
        sel<=2;
        #10
        in0<=4'b0111;
        in1<=4'b1010;
        in2<=4'b1010;
        in3<=4'b1010;
        sel<=0;
        #10
        in0<=8'b01010101;
        in1<=8'b01111101;
        in2<=8'b01110111;
        in3<=8'b01110100;
        sel<=3;
        #10
        in0<=16'b0101010111110000;
        in1<=16'b0101010111110010;
        in2<=16'b0101011111110000;
        in3<=16'b0101110111110000;
        sel<=0;
        #10
        in0<=8'b01011101;
        in1<=8'b01111101;
        in2<=8'b01100111;
        in3<=8'b10110100;
        sel<=1;
        #10
        in0<=16'b0101110111110000;
        in1<=16'b1101010111110010;
        in2<=16'b0101011111111000;
        in3<=16'b0101110100110000;
        sel<=2;
        #10
        in0<=16'b0000000000000000;
        in1<=16'b0000000000000000;
        in2<=16'b0000000000000000;
        in3<=16'b0000000000000000;
        sel<=0;
        #10
        in0<=16'b1111111111111111;
        in1<=16'b1111111111111111;
        in2<=16'b1111111111111111;
        in3<=16'b1111111111111111;
        sel<=3;
        $finish;
    end   
    
    
endmodule
